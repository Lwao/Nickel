library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mux4x1 is
	port(
		
		);
end mux4x1;

architecture proc_of_mux4x1 of mux4x1 is

begin

end proc_of_mux4x1;